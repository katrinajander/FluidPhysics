`default_nettype none

module collision (input wire clk_in,
                input wire rst_in,
                output logic done_colliding);

    // collide everything in BRAM
    // set done_colliding to 1 when done

endmodule

`default_nettype wire