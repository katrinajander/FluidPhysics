`default_nettype none

module streaming();
    // stream everything in BRAM
    // output 1 when done
endmodule

`default_nettype wire