`timescale 1ns / 1ps
`default_nettype none

module top_level
  (
    input wire          clk_100mhz,
    output logic [15:0] led,
    input wire [15:0]   sw,
    input wire [3:0]    btn,
    output logic [2:0] rgb0, //rgb led
    output logic [2:0] rgb1, //rgb led
    output logic [2:0] hdmi_tx_p, //hdmi output signals (positives) (blue, green, red)
    output logic [2:0] hdmi_tx_n, //hdmi output signals (negatives) (blue, green, red)
    output logic hdmi_clk_p, hdmi_clk_n //differential hdmi clock
   );

  // shut up those RGBs
  assign led = sw;
  assign rgb0 = 0;
  assign rgb1 = 0;

  ///////////////////////// BRAM Instantiation for Lattice

  localparam BRAM_DEPTH = 31570; // Comes from (1280/5)*(720/5) = 205*154 = 31570
                                // actual BRAM made with the GUI is 32768
  localparam BRAM_WIDTH = 8; // Lattice densities are 8 bits
  localparam BRAM_SIZE = $clog2(BRAM_DEPTH);
  logic [8:0][BRAM_SIZE-1:0] addra;
  logic [BRAM_SIZE-1:0] addrb;
  logic [8:0][7:0] lbm_bram_data_read;
  logic [8:0][7:0] lbm_bram_data_write;
  logic lbm_write_enable;
  logic sys_rst;

  //HDMI/video registers
  logic [8:0][7:0] hdmi_read_data;
  always_comb begin
    sys_rst = btn[0];
  end

  //              0        1      2         3       4         5       6        7       8
  // BRAM order: center, north, northeast, east, southeast, south, southwest, west, northwest
  // port A for LBM
  // port B for HDMI
  generate
    genvar i;
    for (i=0; i<9; i=i+1)begin
      //this needs to be named blah. don't change it
       blah lattice_ram (
        .addra(addra[i]), // LBM side addressing
        .clka(clk_buf),
        .dina(lbm_bram_data_write[i]), // from LBM module
        .douta(lbm_bram_data_read[i]), // from LBM module
        .ena(1'b1),
        .wea(lbm_write_enable),
        .addrb(addrb),
        .clkb(clk_pixel), //clock for reading for HDMI
        .dinb(), //no data in from HDMI (empty)
        .doutb(hdmi_read_data[i]), //data to get passed along (through calculation) to HDMI
        .enb(1'b1),
        .web(1'b0) //no writing on this side
      );
    end
  endgenerate

  lbm lbm_state_machine (.clk_in(clk_buf),
                .rst_in(sys_rst),
                .bram_data_in(lbm_bram_data_read),
                .sw_in(sw),
                .btn_in(btn[2]),
                .addr_out(addra),
                .bram_data_out(lbm_bram_data_write),
                .valid_data_out(lbm_write_enable));
 
  logic clk_pixel, clk_5x; //clock lines
  logic locked; //locked signal (we'll leave unused but still hook it up)

  logic clk_buf;
  
  BUFG clk_buffer (.I(clk_100mhz), .O(clk_buf));

  //clock manager...creates 74.25 Hz and 5 times 74.25 MHz for pixel and TMDS
  hdmi_clk_wiz_720p mhdmicw (
      .reset(0),
      .locked(locked),
      .clk_ref(clk_buf),
      .clk_pixel(clk_pixel),
      .clk_tmds(clk_5x));
 
  logic [10:0] hcount; //hcount of system
  logic [9:0] vcount; //vcount of system
  logic hor_sync; //horizontal sync signal
  logic vert_sync; //vertical sync signal
  logic active_draw; //ative draw! 1 when in drawing region.0 in blanking/sync
  logic new_frame; //one cycle active indicator of new frame of info!
  logic [5:0] frame_count; //0 to 59 then rollover frame counter

  //pipelining the sync signals with how long bram + logic for pixel generation takes
  localparam PIXEL_LOGIC_DELAY = 2;
  logic hor_sync_pipe [PIXEL_LOGIC_DELAY-1:0];
  logic vert_sync_pipe [PIXEL_LOGIC_DELAY-1:0];
  logic active_draw_pipe [PIXEL_LOGIC_DELAY-1:0];

  always_ff @(posedge clk_pixel) begin
    hor_sync_pipe[0] <= hor_sync;
    vert_sync_pipe[0] <= vert_sync;
    active_draw_pipe[0] <= active_draw;
    for (int i=1; i<PIXEL_LOGIC_DELAY; i = i+1)begin
      hor_sync_pipe[i] <= hor_sync_pipe[i-1];
      vert_sync_pipe[i] <= vert_sync_pipe[i-1];
      active_draw_pipe[i] <= active_draw_pipe[i-1];
    end
  end
 
  //default instantiation so making signals for 720p
  video_sig_gen mvg(
      .pixel_clk_in(clk_pixel),
      .rst_in(sys_rst),
      .hcount_out(hcount),
      .vcount_out(vcount),
      .vs_out(vert_sync),
      .hs_out(hor_sync),
      .ad_out(active_draw),
      .nf_out(new_frame),
      .fc_out(frame_count));

  logic [7:0] red, green, blue; //red green and blue pixel values for output
  logic [7:0] tp_r, tp_g, tp_b; //color values as generated by test_pattern module
  logic [7:0] pg_r, pg_g, pg_b;//color values as generated by pong game(part 2)
  
  //math to convert hcount, vcount value to rgb using lattice data
  pixel_calculator pixels(.pixel_clk_in(clk_pixel),
                          .test_button(btn[1]),
                          .rst_in(sys_rst),
                          .data_in(hdmi_read_data),
                          .hcount_in(hcount),
                          .vcount_in(vcount),
                          .addr_out(addrb),
                          .red_out(red),
                          .green_out(green),
                          .blue_out(blue));
 
  logic [9:0] tmds_10b [0:2]; //output of each TMDS encoder!
  logic tmds_signal [2:0]; //output of each TMDS serializer!
 
  //three tmds_encoders (blue, green, red)
  //note green should have no control signal like red
  //the blue channel DOES carry the two sync signals:
  //  * control_in[0] = horizontal sync signal
  //  * control_in[1] = vertical sync signal
 
  tmds_encoder tmds_red(
      .clk_in(clk_pixel),
      .rst_in(sys_rst),
      .data_in(red),
      .control_in(2'b0),
      .ve_in(active_draw_pipe[PIXEL_LOGIC_DELAY-1]),
      .tmds_out(tmds_10b[2]));

  tmds_encoder tmds_green(
      .clk_in(clk_pixel),
      .rst_in(sys_rst),
      .data_in(green),
      .control_in(2'b0),
      .ve_in(active_draw_pipe[PIXEL_LOGIC_DELAY-1]),
      .tmds_out(tmds_10b[1]));

  tmds_encoder tmds_blue(
      .clk_in(clk_pixel),
      .rst_in(sys_rst),
      .data_in(blue),
      .control_in({vert_sync_pipe[PIXEL_LOGIC_DELAY-1], hor_sync_pipe[PIXEL_LOGIC_DELAY-1]}),
      .ve_in(active_draw_pipe[PIXEL_LOGIC_DELAY-1]),
      .tmds_out(tmds_10b[0]));
 
  //three tmds_serializers (blue, green, red):
  tmds_serializer red_ser(
      .clk_pixel_in(clk_pixel),
      .clk_5x_in(clk_5x),
      .rst_in(sys_rst),
      .tmds_in(tmds_10b[2]),
      .tmds_out(tmds_signal[2]));

  tmds_serializer green_ser(
      .clk_pixel_in(clk_pixel),
      .clk_5x_in(clk_5x),
      .rst_in(sys_rst),
      .tmds_in(tmds_10b[1]),
      .tmds_out(tmds_signal[1]));

  tmds_serializer blue_ser(
      .clk_pixel_in(clk_pixel),
      .clk_5x_in(clk_5x),
      .rst_in(sys_rst),
      .tmds_in(tmds_10b[0]),
      .tmds_out(tmds_signal[0]));
 
  //output buffers generating differential signals:
  //three for the r,g,b signals and one that is at the pixel clock rate
  //the HDMI receivers use recover logic coupled with the control signals asserted
  //during blanking and sync periods to synchronize their faster bit clocks off
  //of the slower pixel clock (so they can recover a clock of about 742.5 MHz from
  //the slower 74.25 MHz clock)
  OBUFDS OBUFDS_blue (.I(tmds_signal[0]), .O(hdmi_tx_p[0]), .OB(hdmi_tx_n[0]));
  OBUFDS OBUFDS_green(.I(tmds_signal[1]), .O(hdmi_tx_p[1]), .OB(hdmi_tx_n[1]));
  OBUFDS OBUFDS_red  (.I(tmds_signal[2]), .O(hdmi_tx_p[2]), .OB(hdmi_tx_n[2]));
  OBUFDS OBUFDS_clock(.I(clk_pixel), .O(hdmi_clk_p), .OB(hdmi_clk_n));

endmodule // top_level
`default_nettype wire

